library verilog;
use verilog.vl_types.all;
entity brent_kung_adder_16bit_tb is
end brent_kung_adder_16bit_tb;
